module sqrt #(
    parameter DW = 64 						//��������λ��
)(
    input wire clk,							//ʱ��
    input wire rst_n,						//�͵�ƽ��λ���첽��λͬ���ͷ�

    input wire [DW-1:0] din_i,				//������������
    input wire din_valid_i,					//����������Ч

    output wire busy_o,						//sqrt��Ԫ��æ

    output wire [(DW+(DW%2))/2-1:0] sqrt_o,	//����������
    output wire [DW-2:0] rem_o				//�����������
);
//��������λ��������չ��ż��
localparam din_width = DW + (DW%2);
//��������
localparam iteration_number = din_width/2;
//����������λ��
localparam icnt_width = clogb2(iteration_number);
//�������λ��
localparam sqrt_width = iteration_number;

//������������Ĵ���
reg [din_width-1:0]din_reg;
//����������
reg [icnt_width-1:0]icnt;
//����״̬�Ĵ�����1;�����У�0:�ȴ�
reg sqrt_en;
//��������Ĵ���
reg [sqrt_width-1:0]sqrt_data;
//��������/���������Ĵ���
reg [DW-2:0]rem_data;

//�������2λ+1
wire [DW:0]sqrt_l2a1 = {sqrt_data, 2'b01};
//�����������¸�2λ�ϳ�
wire [DW:0]rem_a2b = {rem_data, din_reg[din_width-1:din_width-2]};
//�Ƚ�
wire rem_cmp = (rem_a2b>=sqrt_l2a1) ? 1'b1 : 1'b0;
//��һ����������
wire [DW-2:0]rem_next = rem_cmp ? (rem_a2b-sqrt_l2a1) : rem_a2b;
//��һ�����ֽ��
wire sqrt_next = rem_cmp;


//״̬����
always @(posedge clk or negedge rst_n) begin
    if (~rst_n) begin
        sqrt_en <= 1'b0;
        icnt <= iteration_number-1;
    end
    else begin
        case (sqrt_en)
            1'b0 : begin//�ȴ���
                if (din_valid_i) begin//������Ч
                    sqrt_en <= 1'b1;
                    icnt <= iteration_number-1;
                    din_reg <= {{(DW%2){1'b0}}, din_i};//����������չ��ż��
                    sqrt_data <= 0;
                    rem_data <= 0;
                end
            end
            1'b1 : begin//������
                icnt <= icnt-1;
                din_reg <= {din_reg[din_width-3:0], 2'b00};
                sqrt_data <= {sqrt_data[sqrt_width-2:0], sqrt_next};
                rem_data <= rem_next;
                if (icnt==0) begin//��������
                    sqrt_en <= 1'b0;
                end
            end
        endcase
    end
end

assign busy_o = sqrt_en;

assign sqrt_o = sqrt_data;
assign rem_o = rem_data;

//����log2
function integer clogb2;
    input integer depth;
        for (clogb2=0; depth>0; clogb2=clogb2+1)
            depth = depth >> 1;
endfunction
endmodule