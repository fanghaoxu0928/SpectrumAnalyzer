module edge_spy(

      input                  clk,
	  input                  rst_n,
      input                  data,
		
      output                 pos_edge,    //������
	  output                 neg_edge,    //�½���  
	  output                 data_edge,  //���ݱ���
		
	  output reg     [1:0]   D      
);

	always @(posedge clk or negedge rst_n)begin
	    if(rst_n == 1'b0)begin
	        D <= 2'b00;
	    end
	    else begin
	        D <= {D[0], data};  	//D[1]��ʾǰһ״̬��D[0]��ʾ��һ״̬�������ݣ� 
	    end
	end
	
//����߼����б��ؼ��

	assign  pos_edge = ~D[1] & D[0];
	assign  neg_edge = D[1] & ~D[0];
	assign  data_edge = pos_edge | neg_edge;
	
endmodule