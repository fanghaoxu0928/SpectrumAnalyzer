module key_filter
#(
parameter CNT_MAX = 20'd999_999 //�������������ֵ
)
(
input wire sys_clk , //ϵͳʱ�� 50MHz
input wire sys_rst_n , //ȫ�ָ�λ
input wire key_in , //���������ź�

output reg key_flag //key_flag Ϊ 1 ʱ��ʾ�������⵽����������
//key_flag Ϊ 0 ʱ��ʾû�м�⵽����������
);

//********************************************************************//
//****************** Parameter and Internal Signal *******************//
//********************************************************************//
//reg define
reg [19:0] cnt_20ms ; //������

//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//

//cnt_20ms:���ʱ�ӵ������ؼ�⵽�ⲿ���������ֵΪ�͵�ƽʱ����������ʼ����
always@(posedge sys_clk or negedge sys_rst_n)
if(sys_rst_n == 1'b0)
cnt_20ms <= 'd0;
else if(key_in == 1'b1)
cnt_20ms <= 'd0;
else if(cnt_20ms == CNT_MAX && key_in == 1'b0)
cnt_20ms <= cnt_20ms;
else
cnt_20ms <= cnt_20ms + 1'b1;

//key_flag:�������� 20ms �����������Ч��־λ
//�� key_flag �� 999_999 ʱ����,ά��һ��ʱ�ӵĸߵ�ƽ

always@(posedge sys_clk or negedge sys_rst_n)
if(sys_rst_n == 1'b0)
key_flag <= 1'b0;
else if(cnt_20ms == CNT_MAX - 1'b1)
key_flag <= 1'b1;
else
key_flag <= 1'b0;

endmodule