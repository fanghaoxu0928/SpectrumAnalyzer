module fft_top (
    input           i_aclk,         // ʱ���ź�
    input           i_aresetn,      // �첽��λ������Ч��
    input  [15:0]   i_real_data,    // ����ʵ����8λ��
    input           i_data_valid,   // ����������Ч
    input           i_data_last,    // ��������֡������1024�����һ�����ݣ�
    output [63:0]   o_fft_data,     // FFT������ݣ�48λ��ʵ��24λ+�鲿24λ��
    output          o_fft_valid,    // FFT�����Ч
    output          o_fft_last,     // FFT���֡����
    output [23:0]   o_fft_user,     // FFT�û��źţ�ͨ��ΪƵ��������
    output [2:0]    o_alm,          // �澯�ź�
    output          o_stat          // ״̬�ź�
);

// ------------------------------------------------------
// �źŸ�ʽת����8λʵ�� + 8λ�鲿����0���� 16λAXI4S����
// ------------------------------------------------------
reg [31:0] axi4s_data_tdata;
reg        axi4s_data_tvalid;
reg        axi4s_data_tlast;

always @(posedge i_aclk or negedge i_aresetn) begin
    if (!i_aresetn) begin
        axi4s_data_tdata  <= 32'd0;
        axi4s_data_tvalid <= 1'b0;
        axi4s_data_tlast  <= 1'b0;
    end else begin
        // �鲿��0��ʵ����չ��8λ��������Ϊ8λ��ֱ��ƴ�ӣ�
        axi4s_data_tdata  <= {16'd0, i_real_data};  // [31:16]�鲿=0��[15:0]ʵ��=����
        axi4s_data_tvalid <= i_data_valid;          // ����������Ч�ź�
        axi4s_data_tlast  <= i_data_last;           // ����֡�����ź�
    end
end

// ------------------------------------------------------
// ʵ����1024��FFT IP�ˣ�����IP���ɵ�ģ���޸ģ�
// ------------------------------------------------------
fft u_fft (
    .i_axi4s_data_tdata  (axi4s_data_tdata),   // �������ݣ�16λ���鲿8λ+ʵ��8λ��
    .i_axi4s_data_tvalid (axi4s_data_tvalid),  // ������Ч
    .i_axi4s_data_tlast  (axi4s_data_tlast),   // ����֡����
    .o_axi4s_data_tready (),                   // ���������δʹ�ã�����ʼ�վ�����
    .i_axi4s_cfg_tdata   ( 'd0),               // �������ݣ�Ĭ��0��ʹ��IP��Ĭ�����ã�
    .i_axi4s_cfg_tvalid  (1'b0),               // ������Ч��Ĭ��0������̬���ã�
    .i_aclk              (i_aclk),             // ʱ��
    .o_axi4s_data_tdata  (o_fft_data),         // ������ݣ�48λ���鲿24λ+ʵ��24λ��
    .o_axi4s_data_tvalid (o_fft_valid),        // �����Ч
    .o_axi4s_data_tlast  (o_fft_last),         // ���֡����
    .o_axi4s_data_tuser  (o_fft_user),         // ���������0~1023��
    .o_alm               (o_alm),              // �澯
    .o_stat              (o_stat)              // ״̬
);

endmodule